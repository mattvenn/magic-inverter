magic
tech sky130A
timestamp 1592753818
<< nwell >>
rect 31 -1 57 27
<< ntransistor >>
rect 43 -17 46 -7
<< ptransistor >>
rect 43 6 46 16
<< ndiffusion >>
rect 42 -17 43 -7
rect 46 -17 47 -7
<< pdiffusion >>
rect 42 6 43 16
rect 46 6 48 16
<< ndcontact >>
rect 38 -17 42 -7
rect 47 -17 51 -7
<< pdcontact >>
rect 38 6 42 16
rect 48 6 52 16
<< psubstratepcontact >>
rect 34 -28 38 -24
rect 43 -28 47 -24
rect 51 -28 55 -24
<< nsubstratencontact >>
rect 34 20 38 24
rect 42 20 46 24
rect 50 20 54 24
<< polysilicon >>
rect 43 16 46 19
rect 43 -1 46 6
rect 35 -4 46 -1
rect 43 -7 46 -4
rect 43 -20 46 -17
<< polycont >>
rect 31 -4 35 0
<< metal1 >>
rect 32 20 34 24
rect 38 16 42 24
rect 46 20 50 24
rect 54 20 56 24
rect 48 0 52 6
rect 29 -4 31 0
rect 35 -4 36 -1
rect 48 -4 59 0
rect 48 -7 56 -4
rect 38 -24 42 -17
rect 32 -28 43 -24
rect 47 -28 51 -24
rect 55 -28 57 -24
<< labels >>
rlabel metal1 54 20 56 24 6 vdd!
rlabel metal1 29 -4 29 0 1 in
rlabel metal1 59 -4 59 0 7 out
rlabel metal1 47 -28 51 -24 1 gnd!
<< end >>
