.include NMOS-180nm.lib
.include PMOS-180nm.lib

* SPICE3 file created from inverter.ext - technology: min2

.option scale=0.09u

M1000 out in gnd gnd nfet w=10 l=3
+  ad=50 pd=30 as=50 ps=30
M1001 out in vdd vdd pfet w=10 l=3
+  ad=60 pd=32 as=50 ps=30
C0 out gnd 3.26fF
C1 vdd gnd 4.39fF
Vdd vdd gnd 1.8
Vin in gnd pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00
.control
run
plot in out
.endc
.end

