
* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8
Vreset RESET_B VGND 1.8
* Vd D VGND 1.8

* create pulse
Vclk CLK VGND pulse(0 1.8 1n 50p 50p 1n 2n)

* output goes low
*Vd D VGND pulse(1.8 0 942p 50p 50p 2n 2n)
* output goes high
Vd D VGND pulse(1.8 0 943p 50p 50p 2n 2n)

.tran 10e-12 2e-09 0e-00

.control
run
set color0 = white
set color1 = black
plot Q D CLK
.endc

.end
