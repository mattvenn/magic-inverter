* NGSPICE file created from inverter4.ext - technology: sky130A


* Top level circuit inverter4

X0 Y A VPWR NWELL sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 Y A VGND VSUBS sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.end

