Inverter Simulation
* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

* instantiate the inverter
Xinv Y A VPWR VGND VGND VPWR inverter

.subckt inverter Y A NWELL VSUBS VGND VPWR
* NGSPICE file created from inverter.ext - technology: sky130A


* Top level circuit inverter

X0 Y A VPWR NWELL sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 Y A VGND VSUBS sky130_fd_pr__nfet_01v8 w=650000u l=150000u


.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00

.control
run
plot A Y
.endc

.end
