Inverter Simulation
* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

* instantiate the inverter
Xflop CLK D RESET_B VGND VGND VPWR VPWR Q sky130_fd_sc_hd__dfrtp_1 

