* this file edited to remove everything not in tt lib
.lib "./sky130_fd_pr/models/sky130.lib.spice" tt

* instantiate the inverter
Xinv Y A VPWR VGND VGND VPWR sky130_fd_sc_hd__inv_1

