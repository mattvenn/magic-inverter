.include NMOS-180nm.lib
.include PMOS-180nm.lib

