.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00

.control
run
plot A Y
.endc

.end
