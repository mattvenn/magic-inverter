Vdd vdd gnd 1.8
Vin in gnd pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00
.control
run
plot in out
.endc
.end

