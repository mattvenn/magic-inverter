.include sky130_fd_pr/models/sky130.lib.spice

